`define ROW_ADDR_BIT 17
`define SP_CNT_BIT 10
`define N_ENTRY 2720
`define ADDR_CAM_DATA_WIDTH `ROW_ADDR_BIT
`define COUNT_CAM_DATA_WIDTH `SP_CNT_BIT
`define BANK_BITS 32